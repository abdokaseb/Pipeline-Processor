LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;


package Types is
    type ARRAYOFREGS is array(natural range <>) of std_logic_vector;
end package;